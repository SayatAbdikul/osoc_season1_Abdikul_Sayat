module Branch (
    input pc,
    
    output new_pc
);
    
endmodule